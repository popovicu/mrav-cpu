parameter MRAV_ADDR_WIDTH = 16;
parameter MRAV_DATA_WIDTH = 16;
parameter MRAV_REG_NUM = 16;